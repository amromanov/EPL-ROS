module powerlink_rhub_pdo_recv #(parameter master = 0   //?Y?�N�?�???�N�N� ????N�?�???�?�N??�N�, N�N�?? ?????�?�?�?? ???�?????�N�N?
)(                                                      //??????N??�N? ?�?�??N�??N? ??N� ???�N?N�?�N�?� ???�?? ??N�???�N� ??N� N??�?�?????�
    input rst,                     //??N?????N�N�??????N�?? N??�N�??N?
    input clk,                     //???�??N�????N�?? ???�???�N�?�N�??N�
    input [7:0]node,               //????N? node powerlink, ????N�??N�N�?? ???�???? ?�?�N�?�?�?�N�????N�?????�N�N?
    /*input rm_clk,*/                  //RMI Clock    
    input [1:0]rm_rx,              //RMI Rx
    input rm_crs_dv,               //RMI CRS
    output reg pdo_st              //??N�N�???� ??N�??N�?????� ???�???�N�?�
	 //inout [35:0] control
);

wire rx_rdy;                //??N�N�???� ??N�??N�?????� ??N�?�N�?�?????????? ?�?�??N�?�
wire [7:0]rx_data;          //?"?�????N�?� ???� ??N�?�N�?�?????????? ?�?�??N�?�
wire rx_busy;               //?�?�?�?? N�??????, N�N�?? ?????�N� ethernet ???�???�N�

/*rmii_recv_byte rmii_recv_byte(
	.rst(rst),
	.clk(clk),
	.rmii_clk(rm_clk),
	.fast_eth(1),
	.rm_rx_data(rm_rx),
	.rm_crs_dv(rm_crs_dv),
	.data(rx_data),
	.rdy(rx_rdy),
	.busy(rx_busy)
);*/
rmii_recv_byte_50_MHz rmii_recv_byte (
	.rst(rst),
	.clk(clk),
	.fast_eth(1'b1),
	.rm_rx_data(rm_rx),
	.rm_crs_dv(rm_crs_dv),
	.data(rx_data),
	.rdy(rx_rdy),
	.busy(rx_busy)
);

reg [11:0] state_m;        //??N??�??????N�?? ???????�N� ??N�????N?N�?????? ?�?�??N�?� ???�?? st_idle (12 ?�??N�, N�N�???�N� N�??N�???? ???�N�?�???�N�??N�N? Ethernet ???�???�N� ?�NZ?�?????? N�?�?�???�N�?�)
parameter st_idle = 8;     //C??N?N�??N??????� ???�?????�????N? (???�N? N??????�N?N�???� ??N�?�N�?�?? ???????�N� ???�N�???????? ?�?�??N�?� ????N??�?� ??N�???�???�N??�N�) 

reg [8:0]cmp_data;         //?"?�????N�?�, ????N�??N�N�?� ???�???? N?N�?�??????N�N? ?? ??N�?????????�?�?????? ???�???�N�?�, N�N�???�N� ??????N?N�N?, N�N�?? ?�???? ???�???? ??N�N??�??N�N?. ?�????????N�?� ?? 9 ?�??N�?� ???�???�N�?�?�N�, N�N�?? N?N�???? ?�?�??N� N?N�?�?????????�N�N? ???� ???�????
                           //??.?�. cmp_data=9'd256 ???�???�???�N�?�?�N� '???� ??N�?????�N�N?N�N?'
always @(posedge clk, posedge rst)
    if(rst)
        cmp_data = 9'd256;
    else
    case(state_m)   //?' case ??N??� ???????�N� N????�??N?N??�??N� ???� 1, N�.??. cmp_data ???�????????N�N?N? N�???�N????? ???� N??�?�??N?NZN�?�?? N�?�??N�?� ????N??�?� ??N�??N�?????� N?????N�???�N?N�??N?NZN�?�???? ?�???�N�?�????N? state_m
      default  : cmp_data = 9'd256;     //?'N??� ?�?�??N�N� ???� ??????N??�????N�?� ?????�?� ?? case ???� ??N�?????�N�N?NZN�N?N?
//--------------Ethernet ???�???�N�--------------//
            20 : cmp_data = 9'h88;      //?????? ??N�??N�???????�?� - IP (0x88AB)        
            21 : cmp_data = 9'hAB;          
//--------------Powerlink ???�???�N�-------------//
            22 : begin                           //?????? N??????�N�?�????N?
                    if(master)                   
                        cmp_data = {1'b0,/*rx_data[7],*/8'h03};  //?"?�N? ???�N?N�?�N�?� PReq
                    else
                        cmp_data = {1'b0,/*rx_data[7],*/8'h04};  //?"?�N? N??�?�?????� PRes
                 end     
            23 : begin                           //Node ??N?N�??N�???????� (??N�??N�?�??????N??�???? N?N?N�N�????N?N�???�)
                    if(!master)                   
                        cmp_data = 9'd256;       //?"?�N? ???�N?N�?�N�?� ???� ??N�?????�N�N??�N�N?N?
                    else
                        cmp_data = 9'd256;  //?"?�N? N??�?�?????� ??N?N�??N�?????????? ?????�?�?�?? ?�N�N�N? ????N�?�???�?�?�????N�?? node
                 end 
            24 : begin                           //Node ??N�???�?????????� (N?N?N�N�????N?N�???� ????N�??N�????N? ????N??�?�?�??)
                    if(!master)                   
                        cmp_data = 9'd256;  //?"?�N? ???�N?N�?�N�?� N?N�?? ?????�?�?�?? ?�N�N�N? ???????�N� N�?�?�?�N�????N�N??�???????? N??�?�?????�
                    else
                        cmp_data = 9'd256;       //?"?�N? N??�?�?????� ???� ??N�?????�N�N??�N�N?N?
                 end   
         endcase

///reg [8:0]cmp_data2; 		 
//always @(posedge clk, posedge rst)
//    if(rst)
//        cmp_data2 = 9'd256;
//    else
//    case(state_m)   //?' case ??N??� ???????�N� N????�??N?N??�??N� ???� 1, N�.??. cmp_data ???�????????N�N?N? N�???�N????? ???� N??�?�??N?NZN�?�?? N�?�??N�?� ????N??�?� ??N�??N�?????� N?????N�???�N?N�??N?NZN�?�???? ?�???�N�?�????N? state_m
//      default  : cmp_data2 = 9'd256;     //?'N??� ?�?�??N�N� ???� ??????N??�????N�?� ?????�?� ?? case ???� ??N�?????�N�N?NZN�N?N?
////--------------Ethernet ???�???�N�--------------//         
////--------------Powerlink ???�???�N�-------------//
//            22 : begin                           //?????? N??????�N�?�????N?
//                    if(master)                   
//                        cmp_data2 = {1'b0,/*rx_data[7],*/8'h05};  //?"?�N? ???�N?N�?�N�?� PReq
//                    else
//                        cmp_data2 = {1'b0,/*rx_data[7],*/8'h06};  //?"?�N? N??�?�?????� PRes
//                 end        
//         endcase		 
		 
		 
		 
		 
		 
    parameter  last_head = 25; //???????�N� ????N??�?�?????�???? ?�???�?�???�??N�N??�???????? ?�?�??N�?� ???�???�N�?�. ???� ??N?N??????? N??�N?N�?�?? 
                               //??N�?�N�?�?? ???� 1 ?�???�N?N??� ????N??�?�?????�???? ?�?�??N�?�, ????N�??N�N�?? ???�N? ????N�?�N�?�N?N??�N�,
                               //N�N�???�N� N�??N�???? ??N??� ???�N�?�?�??N�?�N�N?
    
    reg fault;      //???�N??�?�?�???�N? ???�N�?�???�?????�N?, ???????�?�N�???�NZN�?�N?, N�N�?? ??N�?????????�?�??N�?? ?? ???�??????N�?? ???????�??N� ???�???�N� ???� ????N�N�?�??N�?�??
    reg head;       //???�N??�?�?�???�N? ???�N�?�???�?????�N?, ???????�?�N�???�NZN�?�N?, N�N�?? ???�N?N? ?�?�?????�???????? N?N????�N????? ??N�????N?N�    

	always @(posedge clk or posedge rst)
		if(rst)
			begin
				state_m <= st_idle; 
                fault <= 0;
                pdo_st <= 0;
                head <= 0;
			end	else 
			begin		
              if(pdo_st)              //????N�?? N??�N�??N? N????????�?�?� pdo_st
                  pdo_st <= 0;  
			   if(rx_busy)            //?�N??�?? ??N�?????????�?�N�N?N? ???�???�N�
			   begin
                   if(rx_rdy&(~head))
                   begin
                      state_m <= state_m + 1;
                      if(~((cmp_data[7:0]==rx_data)||cmp_data[8]))  //?�N??�?? ?�?�??N� ???�???? ??N�?????�N�N?N�N? ?? ???? ???� N�?�???�?? N�????N? ?�???�N�?�????NZ, ????N�??N�????N? ?�N� ???? ?????�?�?�?? ?�N�?� ?�N� ?�N�N�N? N�?�???�??
						//if(!((cmp_data2[7:0] == rx_data) || (cmp_data2 == 9'd256)))  
						  fault <= 1;                                 //???�N�????N�N??�?? ???�????N�?? ???�???�N�, ???�?? ?�??N�N�??
                      if(state_m==last_head)     //?�N??�?? ??N�????N?N� ????N??�?�???????? ?�?�??N� ?�?�?????�???????�, N�??
                        head <= 1;               //??N�N?N�?�???�N??�?? N�?�?�?? head ?? ?�???�N?N??� ????N�?�???? ???� ??N�?????�N�N??�??
                   end
               end else
                   begin
                       if(state_m!=st_idle)                 //?�N??�?? N�???�N????? N�N�?? ?�?�???�N�N????�N?N? ??N�??N'?? ???�???�N�?�
                       begin
                         if(~fault)                         //?�N??�?? ???�???�N� ?�N�?� ??N�????N?N� ?�?�?� ??N????�????
                            pdo_st <= 1;                    //N�?? ??N�N?N�?�???�N??�?? N?N�N�???� pdo_st    
                       end
                       //?'???�??N�?�N�?�?�?? N??�N??�?�?�??N�?� ???�N�?�???�????N�?� ?? ???�N�?�?�N???N�?� N???N?N�??N?????N?
                       state_m <= st_idle;
                       fault   <= 0;
                       head <= 0;
                   end
            end





/*pdo_recv_ila YourInstanceName (
    .CONTROL(control), // INOUT BUS [35:0]
    .CLK(clk), // IN
    .TRIG0(cmp_data), // IN BUS [8:0]
    .TRIG1(rx_data), // IN BUS [7:0]
    .TRIG2(state_m), // IN BUS [11:0]
    .TRIG3(fault), // IN BUS [0:0]
    .TRIG4(head) // IN BUS [0:0]
); */




endmodule
