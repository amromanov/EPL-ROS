module rmii_recv_byte_50_MHz(
    input rst,                  //Асинхронный сброс
    input clk,                  //Тактовый генератор 50 МГц
    input fast_eth,             //Скорость передачи 0 - 10 Мбит/с, 1 - 100 МБит/с  
    input [1:0]rm_rx_data,      //Данные, полученные от phy
    input rm_crs_dv,            //Сигнал phy о наличия принимаемого пакета 
    output reg [7:0]data,       //Данные, полученные по сети
    output reg rdy,             //Сигнал готовности очередного
    output reg busy             //Осуществляется прием пакета (поднимается после идентификации приамбулы и опускает после оконгчания передачи) 
);

//Стробирование входных сигналов
reg [1:0]s_rm_rx_data;
reg s_rm_crs_dv;

always @(posedge rst, posedge clk)
    if(rst)
        {s_rm_rx_data,s_rm_crs_dv} <= 0;
    else
        {s_rm_rx_data,s_rm_crs_dv} <= {rm_rx_data,rm_crs_dv};

reg [4:0]wait_cnt;      //Счетчик ожидания для передачи со скоростью 10 Мбит/c     
reg [7:0]rx_data;       //Регистр принятых данных

reg [1:0]stop;          //Регистр, используемый для грязного хака, позволяющего получить еще один байт после того, как CRS_DV примет низкий уровень в 10 МБитной сети, т.к. почему-то там этот сигнал опускается всегда на 1 байт раньше чем надо 

//Основная логика приёма
always @(posedge rst, posedge clk)
    if(rst)
    begin
        data <= 0;
        rx_data <= 0;
        wait_cnt <= 0;
        rdy <= 0;
        busy <= 0;
        stop <= 0;
    end else
        begin
            if(rdy)         //Автоматически сбрасываем сигнал rdy, чтобы он не длился более 1 такта
                rdy <= 0;
            if(wait_cnt==0)
            begin
                if(!busy)
                begin
                    stop <= 0;              //Снимаем флаг до прихода пакета
                    if(s_rm_crs_dv)         //Если на выходе phy валидные данные
                    begin         
                        if(rx_data==8'hD5)  //Если обнаружили конец преамбулы
                        begin
                            busy <= 1;      //Выставляем сигнал принятия пакета
                            rx_data <= {s_rm_rx_data,6'b11_0000};       //Сохраняем новые данные в rx_data вместе с будующим признаком принятия 1 байта (см. биты 11, которые выдвинутся из регистра}            
                        end else                    
                            rx_data <= {s_rm_rx_data,rx_data[7:2]};     //Пишем кольцом новые данные пока не увидим конец приамбулы 
                        if(!fast_eth)       //В случае 10 Мбитного eth запускаем сторожевой таймер
                            wait_cnt <=9; 
                    end else
                        rx_data <= 0;   //Обнуляем rx_data, чтобы быть уверенными, что сиганл валидности не прерывался
                end else
                    begin
                        if(s_rm_crs_dv|stop[0])            //Если идут валидные байты или принимается последний байт в 10МБитной сети
                        begin
                            if(rx_data[1:0]==2'b11)     //Если принят целый байт
                            begin
                                data <= {s_rm_rx_data,rx_data[7:2]};    //Выводим результат на выход модуля с учетом двух последних принятых бит
                                rx_data <= 8'b11_00_0000;               //Перезагружаем rx_data будующим признаком принятия целого бита
                                if(stop[0])                             //Если принимается последний байт и он уже принят целиком выставляем признак возможности окончить приём пакета
                                    stop <= 2'b10;
                                rdy <= 1;                               //Формируем на выход сигна rdy
                            end else
                                rx_data <= {s_rm_rx_data,rx_data[7:2]}; //В противном случае просто вдвигаем новые 2 бита в rx_data
                            if(!fast_eth)       //В случае 10 Мбитного eth запускаем сторожевой таймер
                                wait_cnt <=9;
                        end else
                            begin       //Если прервался сигнал валидности, то считаем, что пакет принят 
                               if(fast_eth|stop[1])     //Если используется 100 Мбитная сеть или последний байт в 10МБитной сети уже принят
                               begin                    //Оканчиваем приём пакета
                                    stop <= 0;  
                                    busy <= 0;
                                    rx_data <= 0;
                               end else stop <= 2'b01;  //Иначе переходим в режим приёма последнего байта в 10Мбитной сети
                            end
                    end    
            end else
                wait_cnt <= wait_cnt - 1;                               //Уменьщаем счетчик
        end

endmodule
